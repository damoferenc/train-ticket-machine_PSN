--componente necesare pentru componentele sistemului  

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MUX_2_LA_1_1_BIT is 
	port (I0, I1, SEL: in STD_LOGIC;  
	Y: out STD_LOGIC);
end entity MUX_2_LA_1_1_BIT; 

architecture ARHITECTURA_MUX_2_LA_1_1_BIT of MUX_2_LA_1_1_BIT is 
begin  Y <= (I1 and SEL) or (I0 and not (SEL)); 
end ARHITECTURA_MUX_2_LA_1_1_BIT;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MUX_4_LA_1_1_BIT is 
	port (I0, I1, I2, I3, S0, S1: in STD_LOGIC;  
	Y: out STD_LOGIC);
end entity MUX_4_LA_1_1_BIT; 

architecture  ARHITECTURA_MUX_4_LA_1_1_BIT of MUX_4_LA_1_1_BIT is
component MUX_2_LA_1_1_BIT
	port (I0, I1, SEL: in STD_LOGIC;  
	Y: out STD_LOGIC); 
end component;
signal A : STD_LOGIC;
signal B : STD_LOGIC;
begin
	C1:	MUX_2_LA_1_1_BIT port map(I0, I1, S0, A) ;
	C2:	MUX_2_LA_1_1_BIT port map(I2, I3, S0, B) ;
	C3:	MUX_2_LA_1_1_BIT port map(A, B, S1, Y) ; 
end ARHITECTURA_MUX_4_LA_1_1_BIT;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MUX_2_LA_1_4_BIT is 
	port (I0, I1: in STD_LOGIC_VECTOR (0 to 3) ;
	SEL: in STD_LOGIC;  
	Y: out STD_LOGIC_VECTOR ( 0 to 3));
end entity MUX_2_LA_1_4_BIT; 

architecture ARHITECTURA_MUX_2_LA_1_4_BIT of MUX_2_LA_1_4_BIT is 
begin 
	Y(0) <= (I1(0) and SEL) or (I0(0) and not (SEL));
	Y(1) <= (I1(1) and SEL) or (I0(1) and not (SEL));
	Y(2) <= (I1(2) and SEL) or (I0(2) and not (SEL));
	Y(3) <= (I1(3) and SEL) or (I0(3) and not (SEL));
end ARHITECTURA_MUX_2_LA_1_4_BIT;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MUX_4_LA_1_4_BIT is 
	port (I0, I1, I2, I3: in STD_LOGIC_VECTOR ( 0 to 3); 
	S0, S1: in STD_LOGIC;  
	Y: out STD_LOGIC_VECTOR (0 to 3));
end entity MUX_4_LA_1_4_BIT; 

architecture  ARHITECTURA_MUX_4_LA_1_4_BIT of MUX_4_LA_1_4_BIT is
component MUX_2_LA_1_4_BIT is 
	port (I0, I1: in STD_LOGIC_VECTOR (0 to 3) ;
	SEL: in STD_LOGIC;  
	Y: out STD_LOGIC_VECTOR ( 0 to 3)); 
end component;
signal A : STD_LOGIC_vector (0 to 3);
signal B : STD_LOGIC_vector (0 to 3);
begin
	C1:	MUX_2_LA_1_4_BIT port map(I0, I1, S0, A) ;
	C2:	MUX_2_LA_1_4_BIT port map(I2, I3, S0, B) ;
	C3:	MUX_2_LA_1_4_BIT port map(A, B, S1, Y) ; 
end ARHITECTURA_MUX_4_LA_1_4_BIT;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity BISTABIL_D is
	port(D, CLK : in STD_LOGIC;
	Q, NOTQ : out STD_LOGIC);
end BISTABIL_D;

architecture ARHITECTURA_BISTABIL_D of BISTABIL_D is
begin
	process(CLK)
		variable TMP: std_logic;
		begin
			if(CLK='1' and CLK'EVENT) then
				TMP := D;
			end if;
		Q<=TMP;
		NOTQ <=not TMP;
	end PROCESS;
end ARHITECTURA_BISTABIL_D;

library ieee;
use ieee. std_logic_1164.all;
 
entity BISTABIL_JK is
port( J,K,CLOCK: in std_logic;
Q, NOTQ: out std_logic);
end BISTABIL_JK;
 
architecture ARHITECTURA_BISTABIL_JK of BISTABIL_JK is
begin
	process(CLOCK)
	variable TMP: std_logic;
	begin
		if(CLOCK='1' and CLOCK'EVENT) then
			if(J='0' and K='0')then
				TMP:=TMP;
			elsif(J='1' and K='1')then
				TMP:= not TMP;
			elsif(J='0' and K='1')then
				TMP:='0';
			else
				TMP:='1';
			end if;
		end if;
	Q<=TMP;
	NOTQ <=not TMP;
	end PROCESS;
end ARHITECTURA_BISTABIL_JK;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity BCD_7_SEGMENTE is
port ( B0,B1,B2,B3 : in STD_LOGIC;
	   A,B,C,D,E,F,G : out STD_LOGIC);
end BCD_7_SEGMENTE;
 
architecture ARHITECTURA_BCD_7_SEGMENTE of BCD_7_SEGMENTE is
begin
A <= B0 OR B2 OR (B1 AND B3) OR (NOT B1 AND NOT B3);
B <= (NOT B1) OR (NOT B2 AND NOT B3) OR (B2 AND B3);
C <= B1 OR NOT B2 OR B3;
D <= (NOT B1 AND NOT B3) OR (B2 AND NOT B3) OR (B1 AND NOT B2 AND B3) OR (NOT B1 AND B2) OR B0;
E <= (NOT B1 AND NOT B3) OR (B2 AND NOT B3);
F <= B0 OR (NOT B2 AND NOT B3) OR (B1 AND NOT B2) OR (B1 AND NOT B3);
G <= B0 OR (B1 AND NOT B2) OR ( NOT B1 AND B2) OR (B2 AND NOT B3);
end ARHITECTURA_BCD_7_SEGMENTE;	 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity REGISTRU_BCD_8_BIT is
	port(AU, AZ: IN STD_LOGIC_VECTOR(0 TO 3);
	CLK,RESET : IN STD_LOGIC;
	SU, SZ : OUT STD_LOGIC_VECTOR(0 TO 3));
end REGISTRU_BCD_8_BIT;

architecture ARHITECTURA_REGISTRU_BCD_8_BIT of REGISTRU_BCD_8_BIT is
begin
	process(CLK,RESET)
	variable TMPU,TMPZ : std_logic_vector(0 to 3);
	begin
		IF RESET='1' THEN 
			TMPU:="0000" ;
			TMPZ:="0000" ;
		ELSif(CLK = '1' AND CLK'EVENT)	then
			TMPU := AU;
			TMPZ := AZ;
		end if;
		SU <= TMPU;
		SZ <= TMPZ;
	end process;
end ARHITECTURA_REGISTRU_BCD_8_BIT;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity CODIFICATOR is
port ( I50, I20, I10, I5, I2, I1 : in STD_LOGIC;
	   Z0,Z1,Z2,Z3,U0,U1,U2,U3 : out STD_LOGIC);
end CODIFICATOR;
 
architecture ARHITECTURA_CODIFICATOR of CODIFICATOR is
begin
Z3 <= '0';
Z2 <= I50;
Z1 <= I20;
Z0 <= I50 OR I10;
U3 <= '0';
U2 <= I5;
U1 <= I2; 
U0 <= I5 OR I1;
end ARHITECTURA_CODIFICATOR;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity SUMATOR_BCD is
	port(A_U, A_Z, B_U, B_Z : IN STD_LOGIC_VECTOR(0 to 3);
	S_U, S_Z : OUT STD_LOGIC_VECTOR(0 to 3));
end SUMATOR_BCD;

architecture ARHITECTURA_SUMATOR_BCD of SUMATOR_BCD is
begin 
	process(A_Z,A_U,B_Z,B_U)
	variable TU, TZ : std_logic_vector(0 to 3);
	variable COUT : STD_LOGIC;
	begin
		TU := A_U + B_U;
		if(TU > 9 ) then 
			COUT := '1'; 
			TU := TU - 10;
		else
			COUT := '0';
		end if	;
		TZ := A_Z + B_Z+ COUT;
		S_U <= TU;
		S_Z <= TZ;
	end process;
end ARHITECTURA_SUMATOR_BCD;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity NUMARATOR_BCD is 
   port( CLK, MODE: in std_logic; 
   DU, DZ: in std_logic_vector(0 to 3);
 	 RESET, LOAD: in std_logic;
 	 QU, QZ: out std_logic_vector(0 to 3));
end NUMARATOR_BCD;
 
architecture ARHITECTURA_NUMARATOR_BCD of NUMARATOR_BCD is
begin   
	process(CLK,RESET)
	variable TU, TZ: std_logic_vector(0 to 3);
   	begin
      	if RESET='1' then
         	TU := "0000"; 
		 	TZ := "0000";
	  	elsif LOAD='1' and CLK = '1' AND CLK'EVENT then
		 	TU := DU;
		 	TZ := DZ;
      	elsif CLK= '1' and CLK'EVENT and MODE = '1' then
            if TU="1001" then
			   	if TZ="1001" then
				   	TZ:="1001" ;
				   	TU:="1001";
			   	else
				   TZ:= TZ + 1;
				   TU:="0000";
				end if;
			else
				TU := TU+1;
			end if;
	  	elsif (CLK='1' and CLK'EVENT and MODE = '0') then
		   	if TU="0000" then
				if TZ = "0000" then
				   	TU := "0000";
					TZ := "0000";
			   	else
				   TZ := TZ-1 ;
				   TU := "1001";
				end if;
			else
				TU := TU-1;
			end if;
		end if;
		QZ <= TZ;
   		QU <= TU;
   	end process;
end ARHITECTURA_NUMARATOR_BCD;

--componentele sistemului

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MEMORATOR_DE_DISTANTA is
	port(MODE, DIST, INIT, RESET : in std_logic  ;
	DIST_U, DIST_Z : out std_logic_vector(0 to 3));
end MEMORATOR_DE_DISTANTA;

architecture ARHITECTURA_MEMORATOR_DE_DISTANTA of MEMORATOR_DE_DISTANTA is
component NUMARATOR_BCD is 
   port( CLK, MODE: in std_logic; 
   DU, DZ: in std_logic_vector(0 to 3);
 	 RESET, LOAD: in std_logic;
 	 QU, QZ: out std_logic_vector(0 to 3));
end component; 
signal A : STD_LOGIC;
begin
	C1: NUMARATOR_BCD port map(DIST , MODE, "0000", "0000", A, '0', DIST_U, DIST_Z);
	C2: A <= INIT OR RESET;
end ARHITECTURA_MEMORATOR_DE_DISTANTA;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity CALCULATOR_DE_PRET is
	port(DIST_U, DIST_Z : in std_logic_vector(0 to 3);
	PRET_U, PRET_Z : out std_logic_vector (0 to 3));
end CALCULATOR_DE_PRET;

architecture ARHITECTURA_CALCULATOR_DE_PRET of CALCULATOR_DE_PRET is
begin
	PRET_U <= DIST_U;
	PRET_Z <= DIST_Z;
end ARHITECTURA_CALCULATOR_DE_PRET;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity AFISOR_DE_PRET is
	port(PRET_U, PRET_Z : in std_logic_vector(0 to 3);
	SEGMENT_U, SEGMENT_Z : out std_logic_vector(0 to 6));
end AFISOR_DE_PRET;

architecture ARHITECTURA_AFISOR_DE_PRET of AFISOR_DE_PRET is
component BCD_7_SEGMENTE is
port ( B0,B1,B2,B3 : in STD_LOGIC;
	   A,B,C,D,E,F,G : out STD_LOGIC);
end component;
begin
	C1: BCD_7_SEGMENTE port map(PRET_U(0),PRET_U(1),PRET_U(2),PRET_U(3),SEGMENT_U(0),
	SEGMENT_U(1),SEGMENT_U(2),SEGMENT_U(3),SEGMENT_U(4),SEGMENT_U(5),SEGMENT_U(6));
	C2: BCD_7_SEGMENTE port map(PRET_z(0),PRET_z(1),PRET_z(2),PRET_z(3),SEGMENT_z(0),
	SEGMENT_z(1),SEGMENT_z(2),SEGMENT_z(3),SEGMENT_z(4),SEGMENT_z(5),SEGMENT_z(6));	 
end ARHITECTURA_AFISOR_DE_PRET;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity NUMARATOR_DE_BILETE is
	port(DECR, INIT : in STD_LOGIC;
	NUMAR_BILETE : in STD_LOGIC_VECTOR(0 to 3);
	NDB : out STD_LOGIC);
end NUMARATOR_DE_BILETE;

architecture ARHITECTURA_NUMARATOR_DE_BILETE of NUMARATOR_DE_BILETE is
component NUMARATOR_BCD is 
   port( CLK, MODE: in std_logic; 
   DU, DZ: in std_logic_vector(0 to 3);
 	 RESET, LOAD: in std_logic;
 	 QU, QZ: out std_logic_vector(0 to 3));
end component;
SIGNAL S : STD_LOGIC_VECTOR(0 TO 3); 
SIGNAL CLK : STD_LOGIC;
BEGIN
	C1 : NUMARATOR_BCD PORT MAP(CLK,'0', NUMAR_BILETE, "0000", '0', INIT,S);
	C2 : NDB <= S(0) OR S(1) OR S(2) OR S(3);
	C3 : CLK <= DECR OR INIT;
END ARHITECTURA_NUMARATOR_DE_BILETE; 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity COMANDA_PRINTER is
	port(TB, CLK : in STD_LOGIC;
	I2, DECR, PRINTER : out STD_LOGIC);
end COMANDA_PRINTER;

architecture ARHITECTURA_COMANDA_PRINTER of COMANDA_PRINTER is
component BISTABIL_D is
	port(D, CLK : in STD_LOGIC;
	Q, NOTQ : out STD_LOGIC);
end component; 
signal S : STD_LOGIC;
begin
	C1: BISTABIL_D port map(TB, CLK,S );
	I2 <= S;
	DECR <= S;
	PRINTER <= S;
end ARHITECTURA_COMANDA_PRINTER;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY UNITATEA_DE_COMANDA IS
	PORT(I1, START, STOP, CPR, CR, IMP, NDB, I2, CLK, INIT : IN STD_LOGIC;
	SCP, ECR, RBI, R, ELB, EIR, TB : OUT STD_LOGIC);
END UNITATEA_DE_COMANDA;

ARCHITECTURE ARHITECTURA_UNITATEA_DE_COMANDA OF UNITATEA_DE_COMANDA IS
component BISTABIL_D is
	port(D, CLK : in STD_LOGIC;
	Q, NOTQ : out STD_LOGIC);
end component;
COMPONENT MUX_2_LA_1_1_BIT is 
	port (I0, I1, SEL: in STD_LOGIC;  
	Y: out STD_LOGIC);
end COMPONENT;
SIGNAL D0,D1,D2,D3,Q0,Q1,Q2,Q3, NOTQ0, NOTQ1, NOTQ2, NOTQ3, S1, S2, S3, S0 : STD_LOGIC;
BEGIN
	C1 : S3 <= ( Q3 AND Q2 AND NOT Q0) OR(NOT Q2 AND Q1 AND Q0) OR (Q2 AND NOT Q1) OR (NOT Q1 AND NOT Q0)
	OR (NOT NDB AND NOT Q1) OR (NOT I1 AND Q3 AND Q0);
	C2 : S2 <= (Q3 AND NOT Q2 AND NOT Q1) OR (NOT Q3 AND Q0) OR (Q2 AND Q1) OR (STOP AND Q1 AND Q0);
	C3 : S1 <= (Q2 AND NOT Q0) OR (NOT Q3 AND NOT Q2) OR (Q3 AND Q1 AND Q0) OR (STOP AND NOT Q1 AND NOT Q0)
	OR (CR AND Q3 AND Q0) OR (NOT START AND NOT Q3 AND Q1);
	C4 : S0 <= (Q1 AND Q0) OR (NOT Q3 AND Q2 AND Q0) OR (Q3 AND NOT Q1 AND NOT Q0) OR (IMP AND NOT Q1 AND NOT Q0)
	OR (CPR AND Q3 AND NOT Q2) OR (STOP AND Q3 AND Q2 AND Q1) OR (I2 AND NOT Q3 AND Q1);
	C5 : BISTABIL_D PORT MAP(D0, CLK, Q0, NOTQ0); 
	C6 : BISTABIL_D PORT MAP(D1, CLK, Q1, NOTQ1);
	C7 : BISTABIL_D PORT MAP(D2, CLK, Q2, NOTQ2);
	C8 : BISTABIL_D PORT MAP(D3, CLK, Q3, NOTQ3);
	C9 : SCP <= (NOTQ0 AND Q1 AND NOTQ2 AND Q3) or (NOTQ0 AND NOTQ1 AND NOTQ2 AND NOTQ3);
	C10 : ECR <= (NOTQ0 AND NOTQ1 AND NOTQ2 AND Q3) OR (Q0 AND NOTQ1 AND Q2 AND Q3);
	C11 : RBI <= Q0 AND Q1 AND Q2 AND Q3;
	C12 : R <= NOTQ0 AND Q1 AND  Q2 AND NOTQ3;
	C13 : TB <= NOTQ0 AND Q1 AND  Q2 AND NOTQ3;
	C14 : ELB <= NOTQ0 AND Q1 AND Q2 AND Q3;
	C15 : EIR <= Q0 AND Q1 AND NOTQ2 AND Q3;
	C16 : MUX_2_LA_1_1_BIT PORT MAP (S0, '1', INIT, D0);
	C17 : MUX_2_LA_1_1_BIT PORT MAP (S1, '1', INIT, D1);
	C18 : MUX_2_LA_1_1_BIT PORT MAP (S2, '1', INIT, D2);
	C19 : MUX_2_LA_1_1_BIT PORT MAP (S3, '0', INIT, D3);
END ARHITECTURA_UNITATEA_DE_COMANDA;

library IEEE; 
use IEEE.STD_LOGIC_1164.all ;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity CALCULATOR_DE_POSIBILITATE is  
	port(CLOCK, SCP, INIT: in STD_LOGIC;
	REST_U, REST_Z, C1, C2, C5, C10, C20, C50 : IN STD_LOGIC_VECTOR(0 TO 3);
	IMP, CPR: out STD_LOGIC	;
	R1, R2, R5, R10, R20, R50 : OUT STD_LOGIC_VECTOR(0 TO 3));
end CALCULATOR_DE_POSIBILITATE; 
 
architecture ARHITECTURA_CALCULATOR_DE_POSIBILITATE of CALCULATOR_DE_POSIBILITATE is 
type STARE_T is (ST0, ST1, ST2, ST3, ST4, ST5, ST6, ST7); 
signal STARE, NXSTARE: STARE_T; 
SIGNAL RZ, RU, CC1, CC2, CC5, CC10, CC20, CC50, SIGN, RR1, RR2, RR5, RR10, RR20, RR50 : STD_LOGIC_VECTOR(0 TO 3);
begin 
	ACTUALIZEAZ�_STARE: process (INIT, CLOCK) 
	variable VAR_STARE : STARE_T;
	begin   
		if (INIT = '1') then    
			VAR_STARE := ST0;   
		elsif CLOCK'EVENT and CLOCK = '1' then    
			VAR_STARE := NXSTARE;   
		end if; 
		STARE <= VAR_STARE;
	end process ACTUALIZEAZ�_STARE; 
TRANSITIONS: process (STARE, CC1,CC2,CC5,CC10,CC20,CC50, CLOCK)  
begin   
	IMP <= '0'; 
	CPR <= '0'; 
	case STARE is    
		when ST0 => RR1 <= "0000"; RR2 <= "0000"; RR5 <= "0000"; RR10 <= "0000";  RR20 <= "0000"; RR50 <= "0000"; 
			RZ <= REST_Z; RU <= REST_U;
			CC1 <=C1; CC2 <=C2; CC5 <=C5; CC10 <=C10; CC20 <=C20; CC50 <=C50;
			if (SCP = '1') then 
				NXSTARE <= ST1;                    
			else  
				NXSTARE <= ST0;          
			end if;    
		when ST1 =>
			IF (RZ > 4) AND (CC50 > 0) THEN
				RZ <= RZ - 5;
				CC50 <= CC50 - 1;
				RR50 <= RR50 + 1;
				NXSTARE <= ST1;
			ELSE
				NXSTARE <= ST2;	 
			END IF;
		when ST2 => 
			IF (RZ > 1) AND (CC20 > 0) THEN
				RZ <= RZ - 2;
				CC20 <= CC20 - 1;
				RR20 <= RR20 + 1;
				NXSTARE <= ST2;
			ELSE
				NXSTARE <= ST3; 
			END IF;
		when ST3 => 
			IF (RZ > 0) AND (CC10 > 0) THEN
				RZ <= RZ - 1;
				CC10 <= CC10 - 1;
				RR10 <= RR10 + 1;
				NXSTARE <= ST3;
			ELSE
				NXSTARE <= ST4; 
			END IF;
		when ST4 => 
			IF (RU > 4) AND (CC5 > 0) THEN
				RU <= RU - 5;
				CC5 <= CC5 - 1;
				RR5 <= RR5 + 1;
				NXSTARE <= ST4;
			ELSIF (RZ > 0) AND( CC5 > 1) THEN
				RZ <= RZ - 1;
				CC5 <= CC5 - 2;
				RR5 <= RR5 + 2;
				NXSTARE <= ST4;
			ELSE
				NXSTARE <= ST5; 
			END IF;   
		when ST5 => 
			IF (RU > 1) AND (CC2 > 0) THEN
				RU <= RU - 2;
				CC2 <= CC2 - 1;
				RR2 <= RR2 + 1;
				NXSTARE <= ST5;
			ELSIF (RZ > 0) AND (CC2 > 4) THEN
				RZ <= RZ - 1;
				CC2 <= CC2 - 5;
				RR2 <= RR2 + 5;
				NXSTARE <= ST5;
			ELSE
				NXSTARE <= ST6; 
			END IF;    
		when ST6 => 
			IF (RU > 0) AND (CC1 > 0) THEN
				RU <= RU - 1;
				CC1 <= CC1 - 1;	
				RR1 <= RR1 + 1;
				NXSTARE <= ST6;
			ELSIF (RZ > 0) AND (CC1 > 9) THEN
				RZ <= RZ - 1;
				CC1 <= CC1 - 10;
				RR1 <= RR1 + 10;
				NXSTARE <= ST6;
			ELSE
				NXSTARE <= ST7; 
			END IF;    
		when ST7 => 
			IF (RZ > 0) OR (RU > 0) THEN
				IMP <= '1';
				NXSTARE <= ST0;
			ELSE
				CPR <= '1';
				NXSTARE <= ST0;
				R1 <= RR1;
				R2 <= RR2;
				R5 <= RR5;
				R10 <= RR10;
				R20 <= RR20;
				R50 <= RR50;
			END IF;
		end case;  
	end process TRANSITIONS; 
end ARHITECTURA_CALCULATOR_DE_POSIBILITATE;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY CALCULATOR_REST IS
	PORT(ECR, CLK, INIT : IN STD_LOGIC;
	PRET_U, PRET_Z, BANICDF_U, BANICDF_Z : IN STD_LOGIC_VECTOR(0 TO 3);
	CR, EROARE_BANI : OUT STD_LOGIC;
	REST_U, REST_Z : OUT STD_LOGIC_VECTOR (0 TO 3));
END CALCULATOR_REST;

ARCHITECTURE ARHITECTURA_CALCULATOR_REST OF CALCULATOR_REST IS
COMPONENT BISTABIL_JK is
port( J,K,CLOCK: in std_logic;
Q, NOTQ: out std_logic);
end COMPONENT;
component NUMARATOR_BCD is 
   port( CLK, MODE: in std_logic; 
   DU, DZ: in std_logic_vector(0 to 3);
 	 RESET, LOAD: in std_logic;
 	 QU, QZ: out std_logic_vector(0 to 3));
end component;
COMPONENT BISTABIL_D is
	port(D, CLK : in STD_LOGIC;
	Q, NOTQ : out STD_LOGIC);
end COMPONENT;
SIGNAL PL1, PL2, CLK1, CLK2, K1, K2, J1, J2, Q1, Q2, NOTQ1, NOTQ2,R,QD, DELAYED1, DELAYED2, DELAYED3 : STD_LOGIC;
SIGNAL SGU,SGZ,QU, QZ : STD_LOGIC_VECTOR(0 TO 3);
BEGIN
	C1: NUMARATOR_BCD PORT MAP (CLK1, '0', BANICDF_U, BANICDF_Z, R, PL1, SGU, SGZ);
	C2: CLK1 <= CLK AND ECR AND NOT K1;
	C3: NUMARATOR_BCD PORT MAP (CLK2, '0', PRET_U, PRET_Z, INIT, PL2, QU, QZ );
	C5: K1 <= NOT(QU(0) OR QU(1) OR QU(2) OR QU(3) OR QZ(0) OR QZ(1) OR QZ(2) OR QZ(3));
	C6: K2 <= INIT OR DELAYED3;
	C7:	J2 <= ECR;
	C9: BISTABIL_JK PORT MAP (J2, K2, CLK, Q2, NOTQ2);
	C10: PL1 <= NOT(SGU(0) OR SGU(1) OR SGU(2) OR SGU(3) OR SGZ(0) OR SGZ(1) OR SGZ(2) OR SGZ(3));
	C11: PL2 <= ECR AND NOTQ2;
	C12: CR <= K1;
	C13: EROARE_BANI <= ECR AND NOT K1;
	C14: REST_U <= SGU;
	C15: REST_Z <= SGZ;
	C16: CLK2 <= (CLK AND ECR AND NOT QD AND NOT PL1) OR PL2; 
	C17: R <=PL2; 
	C18: BISTABIL_D PORT MAP(PL1,CLK,QD); 
	C19: BISTABIL_D PORT MAP(K1, CLK, DELAYED1);
	C20: BISTABIL_D PORT MAP(DELAYED1, CLK, DELAYED2);
	C21: BISTABIL_D PORT MAP(DELAYED2, CLK, DELAYED3);
END ARHITECTURA_CALCULATOR_REST;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY CODIFICATOR_DE_BANI IS
	PORT(B1,B2,B5,B10,B20,B50 : IN STD_LOGIC;
	BANICDF_U,BANICDF_Z : OUT STD_LOGIC_VECTOR (0 TO 3));
END ENTITY CODIFICATOR_DE_BANI;

ARCHITECTURE ARHITECTURA_CODIFICATOR_DE_BANI OF CODIFICATOR_DE_BANI IS
COMPONENT CODIFICATOR is
port ( I50, I20, I10, I5, I2, I1 : in STD_LOGIC;
	   Z0,Z1,Z2,Z3,U0,U1,U2,U3 : out STD_LOGIC);
end COMPONENT;
BEGIN
	C1: CODIFICATOR PORT MAP (B50, B20, B10, B5, B2, B1, BANICDF_Z(3),BANICDF_Z(2),BANICDF_Z(1),BANICDF_Z(0),
	BANICDF_U(3),BANICDF_U(2),BANICDF_U(1),BANICDF_U(0)); 
END ARHITECTURA_CODIFICATOR_DE_BANI; 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY MEMORATOR_DE_SUMA_INTRODUSA IS
	PORT(BANICDF_U, BANICDF_Z : STD_LOGIC_VECTOR(0 TO 3);
	CLK, INIT, RBI : IN STD_LOGIC;
	SUMA_U, SUMA_Z : OUT STD_LOGIC_VECTOR (0 TO 3));
END MEMORATOR_DE_SUMA_INTRODUSA;

ARCHITECTURE ARHITECTURA_MEMORATOR_DE_SUMA_INTRODUSA OF MEMORATOR_DE_SUMA_INTRODUSA IS
COMPONENT SUMATOR_BCD is
	port(A_U, A_Z, B_U, B_Z : IN STD_LOGIC_VECTOR(0 to 3);
	S_U, S_Z : OUT STD_LOGIC_VECTOR(0 to 3));
end COMPONENT;
COMPONENT REGISTRU_BCD_8_BIT is
	port(AU, AZ: IN STD_LOGIC_VECTOR(0 TO 3);
	CLK,RESET : IN STD_LOGIC;
	SU, SZ : OUT STD_LOGIC_VECTOR(0 TO 3));
end COMPONENT;
SIGNAL SU, SZ, SSU, SSZ : STD_LOGIC_VECTOR (0 TO 3);
SIGNAL RESET : STD_LOGIC;
BEGIN
	C1: SUMATOR_BCD PORT MAP (BANICDF_U, BANICDF_Z, SU, SZ,SSU,SSZ);
	C2 : REGISTRU_BCD_8_BIT PORT MAP(SSU, SSZ,CLK, RESET, SU, SZ);
	C3 : SUMA_U <= SU;
	C4 : SUMA_Z <= SZ; 
	C5 : RESET <= INIT OR RBI;
END ARHITECTURA_MEMORATOR_DE_SUMA_INTRODUSA;

library IEEE; 
use IEEE.STD_LOGIC_1164.all ;

ENTITY MEMORATOR_DE_BANI IS
	PORT(B1, B2, B5, B10, B20, B50, INIT, I1 : IN STD_LOGIC;
	NUM1 ,NUM2, NUM5, NUM10, NUM20, NUM50 : OUT STD_LOGIC_VECTOR(0 TO 3));
END MEMORATOR_DE_BANI;

ARCHITECTURE ARHITECTURA_MEMORATOR_DE_BANI OF MEMORATOR_DE_BANI IS
component NUMARATOR_BCD is 
   port( CLK, MODE: in std_logic; 
   DU, DZ: in std_logic_vector(0 to 3);
 	 RESET, LOAD: in std_logic;
 	 QU, QZ: out std_logic_vector(0 to 3));
end component; 
SIGNAL RESET : STD_LOGIC;
BEGIN
	C1:NUMARATOR_BCD PORT MAP(B1, '1', "0000", "0000", RESET, '0', NUM1 );
	C2:NUMARATOR_BCD PORT MAP(B2, '1', "0000", "0000", RESET, '0', NUM2 );
	C3:NUMARATOR_BCD PORT MAP(B5, '1', "0000", "0000", RESET, '0', NUM5 );
	C4:NUMARATOR_BCD PORT MAP(B10, '1', "0000", "0000", RESET, '0', NUM10 );
	C5:NUMARATOR_BCD PORT MAP(B20, '1', "0000", "0000", RESET, '0', NUM20 );
	C6:NUMARATOR_BCD PORT MAP(B50, '1', "0000", "0000", RESET, '0', NUM50);
	C7:RESET <= INIT OR I1;
END ARHITECTURA_MEMORATOR_DE_BANI;

library IEEE; 
use IEEE.STD_LOGIC_1164.all ;

ENTITY CASA_DE_BANI IS
	PORT(INIT,B1 ,B2 ,B5 ,B10, B20, B50, P1, P2, P5, P10, P20, P50 : IN STD_LOGIC; 
	I1, I2, I5, I10, I20, I50 : IN STD_LOGIC_VECTOR(0 TO 3);
	NUM1 ,NUM2 ,NUM5, NUM10, NUM20, NUM50 : OUT STD_LOGIC_VECTOR (0 TO 3));
END	CASA_DE_BANI;

ARCHITECTURE ARHITECTURA_CASA_DE_BANI OF CASA_DE_BANI IS
component NUMARATOR_BCD is 
   port( CLK, MODE: in std_logic; 
   DU, DZ: in std_logic_vector(0 to 3);
 	 RESET, LOAD: in std_logic;
 	 QU, QZ: out std_logic_vector(0 to 3));
end component; 
component MUX_2_LA_1_1_BIT
	port (I0, I1, SEL: in STD_LOGIC;  
	Y: out STD_LOGIC); 
end component;
SIGNAL CLK1,CLK2,CLK3,CLK4,CLK5,CLK6, M1,M2,M3,M4,M5,M6 : STD_LOGIC; 
BEGIN
	C1:NUMARATOR_BCD PORT MAP(CLK1, M1, I1, "0000", '0',INIT, NUM1 );
	C2:NUMARATOR_BCD PORT MAP(CLK2, M2, I2, "0000", '0',INIT, NUM2 );
	C3:NUMARATOR_BCD PORT MAP(CLK3, M3, I5, "0000", '0',INIT, NUM5 );
	C4:NUMARATOR_BCD PORT MAP(CLK4, M4, I10, "0000", '0',INIT, NUM10 );
	C5:NUMARATOR_BCD PORT MAP(CLK5, M5, I20, "0000", '0',INIT, NUM20 );
	C6:NUMARATOR_BCD PORT MAP(CLK6, M6, I50, "0000", '0',INIT, NUM50); 
	C7:CLK1 <= B1 OR P1 OR INIT; 
	C8:CLK2 <= B2 OR P2 OR INIT;
	C9:CLK3 <= B5 OR P5 OR INIT;
	C10:CLK4 <= B10 OR P10 OR INIT;
	C11:CLK5 <= B20 OR P20 OR INIT;
	C12:CLK6 <= B50 OR P50 OR INIT;
	C13:MUX_2_LA_1_1_BIT PORT MAP('0','1',B1,M1);  
	C14:MUX_2_LA_1_1_BIT PORT MAP('0','1',B2,M2);
	C15:MUX_2_LA_1_1_BIT PORT MAP('0','1',B5,M3);
	C16:MUX_2_LA_1_1_BIT PORT MAP('0','1',B10,M4);
	C17:MUX_2_LA_1_1_BIT PORT MAP('0','1',B20,M5);
	C18:MUX_2_LA_1_1_BIT PORT MAP('0','1',B50,M6);
END ARHITECTURA_CASA_DE_BANI;
			 
library IEEE; 
use IEEE.STD_LOGIC_1164.all ;

ENTITY COMANDA_DE_PLATIRE IS
	PORT(RBI, R, NCLK, INIT : IN STD_LOGIC;
	B1, B2, B5, B10, B20, B50, R1 ,R2, R5, R10, R20, R50 : IN STD_LOGIC_VECTOR (0 TO 3);
	I1,P1 ,P2, P5, P10, P20, P50 : OUT STD_LOGIC);
END COMANDA_DE_PLATIRE;

ARCHITECTURE ARHITECTURA_COMANDA_DE_PLATIRE OF COMANDA_DE_PLATIRE IS
COMPONENT MUX_4_LA_1_4_BIT is 
	port (I0, I1, I2, I3: in STD_LOGIC_VECTOR ( 0 to 3); 
	S0, S1: in STD_LOGIC;  
	Y: out STD_LOGIC_VECTOR (0 to 3));
end  COMPONENT;
COMPONENT BISTABIL_JK is
port( J,K,CLOCK: in std_logic;
Q, NOTQ: out std_logic);
end COMPONENT;
component NUMARATOR_BCD is 
   port( CLK, MODE: in std_logic; 
   DU, DZ: in std_logic_vector(0 to 3);
 	 RESET, LOAD: in std_logic;
 	 QU, QZ: out std_logic_vector(0 to 3));
end component;	
COMPONENT BISTABIL_D is
	port(D, CLK : in STD_LOGIC;
	Q, NOTQ : out STD_LOGIC);
end COMPONENT;
SIGNAL S1, S2, S5, S10, S20, S50, Q1, Q2, Q5, Q10, Q20, Q50 : STD_LOGIC_VECTOR(0 TO 3);
SIGNAL PL,J,K,Q, ECD1, ECD2, ECD5, ECD10, ECD20, ECD50,II,E1,E2,E5,E10,E20,E50,RR, RR1,RR2,RR3,IDELAYED, IFINAL : std_logic;
SIGNAL PP1,PP2,PP5,PP10,PP20,PP50, E1DEL, E2DEL, E5DEL, E10DEL, E20DEL,E50DEL, PLDELAYED, KDELAYED, CLK : STD_LOGIC;
BEGIN
	C1: MUX_4_LA_1_4_BIT PORT MAP("0000",B1,R1, "0000", RBI, R,S1);	
	C2: MUX_4_LA_1_4_BIT PORT MAP("0000",B2,R2, "0000", RBI, R,S2);
	C3: MUX_4_LA_1_4_BIT PORT MAP("0000",B5,R5, "0000", RBI, R,S5);
	C4: MUX_4_LA_1_4_BIT PORT MAP("0000",B10,R10, "0000", RBI, R,S10);
	C5: MUX_4_LA_1_4_BIT PORT MAP("0000",B20,R20, "0000", RBI, R,S20);
	C6: MUX_4_LA_1_4_BIT PORT MAP("0000",B50,R50, "0000", RBI, R,S50);
	C7: NUMARATOR_BCD PORT MAP(ECD1,'0', S1, "0000",INIT,PL, Q1);
	C8: NUMARATOR_BCD PORT MAP(ECD2,'0', S2, "0000",INIT,PL, Q2);
	C9: NUMARATOR_BCD PORT MAP(ECD5,'0', S5, "0000",INIT,PL, Q5);
	C10: NUMARATOR_BCD PORT MAP(ECD10,'0', S10, "0000",INIT,PL, Q10);
	C11: NUMARATOR_BCD PORT MAP(ECD20,'0', S20, "0000",INIT,PL, Q20);
	C12: NUMARATOR_BCD PORT MAP(ECD50,'0', S50, "0000",INIT,PL, Q50);
	C13: BISTABIL_JK PORT MAP(J,K,CLK, Q);
	C14: K <= RBI OR R;
	C15: PL <= Q AND K;
	C16: ECD1 <= (CLK AND K)OR PL;
	C17: ECD2 <= (NOT PP1 AND CLK AND E1DEL) OR PL ;
	C18: ECD5 <= (NOT PP2 AND CLK AND E2DEL AND E1DEL) OR PL;
	C19: ECD10 <= (NOT PP5 AND CLK AND E5DEL AND E2DEL AND E1DEL) OR PL;
	C20: ECD20 <= (NOT PP10 AND CLK AND E10DEL AND E5DEL AND E2DEL AND E1DEL) OR PL;
	C21: ECD50 <= (NOT PP20 AND CLK AND E20DEL AND E10DEL AND E5DEL AND E2DEL AND E1DEL) OR PL;
	C22: J <= INIT OR II;
	C23: II <= E1 AND E2 AND E5 AND E10 AND E20 AND E50;
	C24: PP1 <= ECD1 AND NOT E1DEL AND NOT PL AND NOT PLDELAYED ;
	C25: PP2 <= ECD2 AND NOT E2DEL AND NOT PL AND NOT PLDELAYED	;
	C26: PP5 <= ECD5 AND NOT E5DEL AND NOT PL AND NOT PLDELAYED ;
	C27: PP10 <= ECD10 AND NOT E10DEL AND NOT PL AND NOT PLDELAYED ;	
	C28: PP20 <= ECD20 AND NOT E20DEL AND NOT PL AND NOT PLDELAYED	;
	C29: PP50 <= ECD50 AND NOT E50DEL AND NOT PL AND NOT PLDELAYED	 ;	
	C30: I1<= IDELAYED AND IFINAL AND II AND K; 
	C31: E1 <= NOT(Q1(1)OR Q1(2)OR Q1(3)OR Q1(0));
	C32: E2 <= NOT(Q2(1)OR Q2(2)OR Q2(3)OR Q2(0));
	C33: E5 <= NOT(Q5(1)OR Q5(2)OR Q5(3)OR Q5(0));	
	C34: E10 <= NOT(Q10(1)OR Q10(2)OR Q10(3)OR Q10(0));
	C35: E20 <= NOT(Q20(1)OR Q20(2)OR Q20(3)OR Q20(0));
	C36: E50 <=	NOT(Q50(1)OR Q50(2)OR Q50(3)OR Q50(0));
	C37: BISTABIL_D PORT MAP(II, CLK,IDELAYED);
	C38: BISTABIL_D PORT MAP(IDELAYED, CLK, IFINAL);  
	C39: P1 <= PP1;
	C40: P2 <= PP2;
	C41: P5 <= PP5;
	C42: P10 <= PP10;
	C43: P20 <= PP20;
	C44: P50 <= PP50;
	C45: BISTABIL_D PORT MAP(E1, CLK, E1DEL); 
	C46: BISTABIL_D PORT MAP(E2, CLK, E2DEL);
	C47: BISTABIL_D PORT MAP(E5, CLK, E5DEL);
	C48: BISTABIL_D PORT MAP(E10, CLK, E10DEL);
	C49: BISTABIL_D PORT MAP(E20, CLK, E20DEL);
	C50: BISTABIL_D PORT MAP(E50, CLK, E50DEL);
	C51: BISTABIL_D PORT MAP(PL, CLK, PLDELAYED);
	C52: CLK <= NOT NCLK;
	
END ARHITECTURA_COMANDA_DE_PLATIRE;

--SISTEMUL

library IEEE; 
use IEEE.STD_LOGIC_1164.all ;  

ENTITY AUTOMAT_DE_BILETE IS
	PORT(DIST, MODE, START, STOP, INIT, CLock: IN STD_LOGIC;
	B1, B2, B5, B10, B20, B50: IN STD_LOGIC;
	INN, NR_BILETE : IN STD_LOGIC_VECTOR(0 TO 3);
	RE1, RE2, RE5, RE10, RE20, RE50: OUT STD_LOGIC;
	ANODE : OUT  STD_LOGIC_VECTOR(0 TO 3);
	LED_OUT : OUT STD_LOGIC_VECTOR(0 TO 6); 
	ERROR_BANI, ERROR_BILETE, ERROR_RESTITUIRE, BILET  : OUT STD_LOGIC);
END AUTOMAT_DE_BILETE;

ARCHITECTURE ARHITECTURA_AUTOMAT_DE_BILETE OF AUTOMAT_DE_BILETE IS
COMPONENT MEMORATOR_DE_DISTANTA is
	port(MODE, DIST, INIT, RESET : in std_logic  ;
	DIST_U, DIST_Z : out std_logic_vector(0 to 3));
end COMPONENT;
COMPONENT CALCULATOR_DE_PRET is
	port(DIST_U, DIST_Z : in std_logic_vector(0 to 3);
	PRET_U, PRET_Z : out std_logic_vector (0 to 3));
end COMPONENT;
COMPONENT AFISOR_DE_PRET is
	port(PRET_U, PRET_Z : in std_logic_vector(0 to 3);
	SEGMENT_U, SEGMENT_Z : out std_logic_vector(0 to 6));
end COMPONENT;
COMPONENT NUMARATOR_DE_BILETE is
	port(DECR, INIT : in STD_LOGIC;
	NUMAR_BILETE : in STD_LOGIC_VECTOR(0 to 3);
	NDB : out STD_LOGIC);
end COMPONENT;
COMPONENT COMANDA_PRINTER is
	port(TB, CLK : in STD_LOGIC;
	I2, DECR, PRINTER : out STD_LOGIC);
end COMPONENT;
COMPONENT UNITATEA_DE_COMANDA IS
	PORT(I1, START, STOP, CPR, CR, IMP, NDB, I2, CLK, INIT : IN STD_LOGIC;
	SCP, ECR, RBI, R, ELB, EIR, TB : OUT STD_LOGIC);
END COMPONENT;
COMPONENT CALCULATOR_DE_POSIBILITATE is  
	port(CLOCK, SCP, INIT: in STD_LOGIC;
	REST_U, REST_Z, C1, C2, C5, C10, C20, C50 : IN STD_LOGIC_VECTOR(0 TO 3);
	IMP, CPR: out STD_LOGIC	;
	R1, R2, R5, R10, R20, R50 : OUT STD_LOGIC_VECTOR(0 TO 3));
end COMPONENT;
COMPONENT CALCULATOR_REST IS
	PORT(ECR, CLK, INIT : IN STD_LOGIC;
	PRET_U, PRET_Z, BANICDF_U, BANICDF_Z : IN STD_LOGIC_VECTOR(0 TO 3);
	CR, EROARE_BANI : OUT STD_LOGIC;
	REST_U, REST_Z : OUT STD_LOGIC_VECTOR (0 TO 3));
END COMPONENT;
COMPONENT CODIFICATOR_DE_BANI IS
	PORT(B1,B2,B5,B10,B20,B50 : IN STD_LOGIC;
	BANICDF_U,BANICDF_Z : OUT STD_LOGIC_VECTOR (0 TO 3));
END COMPONENT;
COMPONENT MEMORATOR_DE_SUMA_INTRODUSA IS
	PORT(BANICDF_U, BANICDF_Z : STD_LOGIC_VECTOR(0 TO 3);
	CLK, INIT, RBI : IN STD_LOGIC;
	SUMA_U, SUMA_Z : OUT STD_LOGIC_VECTOR (0 TO 3));
END COMPONENT;
COMPONENT MEMORATOR_DE_BANI IS
	PORT(B1, B2, B5, B10, B20, B50, INIT, I1 : IN STD_LOGIC;
	NUM1 ,NUM2, NUM5, NUM10, NUM20, NUM50 : OUT STD_LOGIC_VECTOR(0 TO 3));
END COMPONENT;
COMPONENT CASA_DE_BANI IS
	PORT(INIT,B1 ,B2 ,B5 ,B10, B20, B50, P1, P2, P5, P10, P20, P50 : IN STD_LOGIC; 
	I1, I2, I5, I10, I20, I50 : IN STD_LOGIC_VECTOR(0 TO 3);
	NUM1 ,NUM2 ,NUM5, NUM10, NUM20, NUM50 : OUT STD_LOGIC_VECTOR (0 TO 3));
END	COMPONENT;
COMPONENT COMANDA_DE_PLATIRE IS
	PORT(RBI, R, NCLK, INIT : IN STD_LOGIC;
	B1, B2, B5, B10, B20, B50, R1 ,R2, R5, R10, R20, R50 : IN STD_LOGIC_VECTOR (0 TO 3);
	I1,P1 ,P2, P5, P10, P20, P50 : OUT STD_LOGIC);
END COMPONENT; 
COMPONENT BISTABIL_D is
	port(D, CLK : in STD_LOGIC;
	Q, NOTQ : out STD_LOGIC);
end COMPONENT;
component DIVIZOR_DE_FRECVENTA		IS
	PORT(CLOCK : IN STD_LOGIC;
	CLK : OUT STD_LOGIC);
END component;
component FPGA_7_SEGMENTE IS
	PORT(CLOCK: IN STD_LOGIC;
	PRET_U, PRET_Z, SUMA_U, SUMA_Z : IN STD_LOGIC_VECTOR(0 TO 6);
	ANODE : OUT  STD_LOGIC_VECTOR(0 TO 3);
	LED_OUT : OUT STD_LOGIC_VECTOR(0 TO 6));
END component;
COMPONENT DEBOUNCE IS
	PORT(D, CLK : IN STD_LOGIC;
	Q : OUT STD_LOGIC);
END COMPONENT;
SIGNAL DECR,NDB,TB,I2,R,I1,RBI,CR,ECR,CPR,SCP,IMP,P1,P2,P5,P10,P20,P50, CLK: STD_LOGIC;
SIGNAL REST_U,REST_Z,DISTANTA_U,DISTANTA_Z,PRET_U,PRET_Z,C1,C2,C5,C10,C20,C50,R1,R2,R5,R10,R20,R50 : STD_LOGIC_VECTOR(0 TO 3);
SIGNAL BANICDF_U,BANICDF_Z,SUMA_U,SUMA_Z,NUM1 ,NUM2, NUM5, NUM10, NUM20, NUM50 : STD_LOGIC_VECTOR(0 TO 3); 
SIGNAL CLKMEMSUM, CLKMEMSUMDELAYED, CPRDELAYED, CPRFINAL, IMPDELAYED, IMPFINAL : STD_LOGIC;
SIGNAL I1DELAYED, RESETCALCULATORREST : STD_LOGIC;
signal clockdivizat, clockdivizat2, clockdivizat3 : STD_LOGIC;
signal SUMAINTR_U, SUMAINTR_Z, COST_U, COST_Z : STD_LOGIC_VECTOR(0 TO 6);
SIGNAL DIST_DEBOUNCED, START_DEBOUNCED,STOP_DEBOUNCED : STD_LOGIC;
SIGNAL IN1, IN2, IN5, IN10, IN20, IN50 : STD_LOGIC_VECTOR(0 TO 3);
BEGIN
	CC1: MEMORATOR_DE_DISTANTA PORT MAP(MODE, DIST_DEBOUNCED,INIT,R,DISTANTA_U,DISTANTA_Z);
	CC2: CALCULATOR_DE_PRET PORT MAP(DISTANTA_U,DISTANTA_Z,PRET_U,PRET_Z);
	CC3: AFISOR_DE_PRET PORT MAP(PRET_U,PRET_Z,COST_U,COST_Z);
	CC4: NUMARATOR_DE_BILETE PORT MAP(DECR, INIT, NR_BILETE,NDB);
	CC5: COMANDA_PRINTER PORT MAP(TB, CLK, I2, DECR, BILET);
	CC6: UNITATEA_DE_COMANDA PORT MAP(I1,START_DEBOUNCED,STOP_DEBOUNCED,CPRFINAL,CR,IMPFINAL,NDB,I2,CLK,INIT,SCP,ECR,RBI,R,ERROR_BILETE,ERROR_RESTITUIRE,TB);
	CC7: CALCULATOR_DE_POSIBILITATE PORT MAP(CLK,SCP,INIT,REST_U,REST_Z,C1,C2,C5,C10,C20,C50,IMP,CPR,R1,R2,R5,R10,R20,R50);
	CC8: CALCULATOR_REST PORT MAP(ECR,CLK,RESETCALCULATORREST,PRET_U,PRET_Z,BANICDF_U,BANICDF_Z,CR,ERROR_BANI,REST_U,REST_Z);
	CC9: CODIFICATOR_DE_BANI PORT MAP(B1,B2,B5,B10,B20,B50,BANICDF_U,BANICDF_Z);
	CC10: MEMORATOR_DE_SUMA_INTRODUSA PORT MAP(BANICDF_U,BANICDF_Z,CLKMEMSUMDELAYED, INIT, RBI,SUMA_U,SUMA_Z);
	CC11: AFISOR_DE_PRET PORT MAP(SUMA_U,SUMA_Z,SUMAINTR_U,SUMAINTR_Z);
	CC12: MEMORATOR_DE_BANI PORT MAP(B1,B2,B5,B10,B20,B50,INIT,I1,NUM1,NUM2,NUM5,NUM10,NUM20,NUM50);
	CC13: CASA_DE_BANI PORT MAP(INIT,B1,B2,B5,B10,B20,B50,P1,P2,P5,P10,P20,P50,IN1,IN2,IN5,IN10,IN20,IN50,C1,C2,C5,C10,C20,C50);
	CC14: COMANDA_DE_PLATIRE PORT MAP(RBI,R,CLockdivizat2,INIT,NUM1,NUM2,NUM5,NUM10,NUM20,NUM50,R1,R2,R5,R10,R20,R50,I1,P1,P2,P5,P10,P20,P50);
	CC15: RE1 <= P1;
	CC16: RE2 <= P2;
	CC17: RE5 <= P5;
	CC18: RE10 <= P10;
	CC19: RE20 <= P20;
	CC20: RE50 <= P50; 
	CC21: CLKMEMSUM <= B1 OR B2 OR B5 OR B10 OR B20 OR B50;	
	CC22: BISTABIL_D PORT MAP(CLKMEMSUM, CLK, CLKMEMSUMDELAYED);
	CC23: BISTABIL_D PORT MAP(CPR, CLK, CPRDELAYED);
	CC24: CPRFINAL <= CPR OR CPRDELAYED;
	CC25: IMPFINAL <= IMPDELAYED OR IMP;
	CC26: BISTABIL_D PORT MAP(IMP, CLK, IMPDELAYED);
	CC27: BISTABIL_D PORT MAP(I1, CLK, I1DELAYED) ;
	CC28: RESETCALCULATORREST <= INIT OR I1;
	cc29: divizor_de_frecventa port map (clock, clk);
	cc30: divizor_de_frecventa port map (clk, clockdivizat);
	cc31: divizor_de_frecventa port map (clockdivizat, clockdivizat2);
	cc32: fpga_7_segmente port map(clk, cost_U, cost_Z, SUMAintr_U, SUMAintr_Z, anode, led_out);
	CC33: DEBOUNCE PORT MAP (START, CLK, START_DEBOUNCED);
	CC34: DEBOUNCE PORT MAP (STOP, CLK, STOP_DEBOUNCED);
	CC35: DEBOUNCE PORT MAP (DIST, CLK, DIST_DEBOUNCED);
	CC36: IN1 <= INN;
	CC37: IN2 <= INN;
	CC38: IN5 <= INN;
	CC39: IN10 <= INN;
	CC40: IN20 <= INN;
	CC41: IN50 <= INN;
	
END ARHITECTURA_AUTOMAT_DE_BILETE;
	





















library IEEE; 
use IEEE.STD_LOGIC_1164.all ;

ENTITY DIVIZOR_DE_FRECVENTA		IS
	PORT(CLOCK : IN STD_LOGIC;
	CLK : OUT STD_LOGIC);
END DIVIZOR_DE_FRECVENTA;

ARCHITECTURE ARHITECTURA_DIVIZOR_DE_FRECVENTA OF DIVIZOR_DE_FRECVENTA IS
COMPONENT BISTABIL_JK is
port( J,K,CLOCK: in std_logic;
Q, NOTQ: out std_logic);
end COMPONENT;
SIGNAL Q1,Q2,Q3,Q4,Q5,Q6: STD_LOGIC;
BEGIN
	C1: BISTABIL_JK PORT MAP('1','1', CLOCK,Q1);
	C2: BISTABIL_JK PORT MAP(Q1,Q1, CLOCK,Q2);
	C3: BISTABIL_JK PORT MAP(Q2,Q2, CLOCK,Q3);
	C4: BISTABIL_JK PORT MAP(Q3,Q3, CLOCK,Q4);
	C5: BISTABIL_JK PORT MAP(Q4,Q4, CLOCK,Q5);
	C6: BISTABIL_JK PORT MAP(Q5,Q5, CLOCK,Q6); 
	C7: CLK <= Q6;
END ARHITECTURA_DIVIZOR_DE_FRECVENTA;

library IEEE; 
use IEEE.STD_LOGIC_1164.all ;

ENTITY DEBOUNCE IS
	PORT(D, CLK : IN STD_LOGIC;
	Q : OUT STD_LOGIC);
END DEBOUNCE;

ARCHITECTURE ARHITECTURA_DEBOUNCE OF DEBOUNCE IS
COMPONENT BISTABIL_D is
	port(D, CLK : in STD_LOGIC;
	Q, NOTQ : out STD_LOGIC);
end COMPONENT;
SIGNAL Q1,Q2,Q3 : STD_LOGIC;
BEGIN
	C1: BISTABIL_D PORT MAP (D, CLK, Q1);
	C2: BISTABIL_D PORT MAP (Q1, CLK, Q2);
	C3: BISTABIL_D PORT MAP (Q2, CLK, Q3);
	C4: Q <= Q1 AND Q2 AND Q3;
END ARHITECTURA_DEBOUNCE;	

library IEEE; 
use IEEE.STD_LOGIC_1164.all ; 
use IEEE.std_logic_unsigned.all;

ENTITY FPGA_7_SEGMENTE IS
	PORT(CLOCK: IN STD_LOGIC;
	PRET_U, PRET_Z, SUMA_U, SUMA_Z : IN STD_LOGIC_VECTOR(0 TO 6);
	ANODE : OUT  STD_LOGIC_VECTOR(0 TO 3);
	LED_OUT : OUT STD_LOGIC_VECTOR(0 TO 6));
END FPGA_7_SEGMENTE;

ARCHITECTURE ARHITECTURA_FPGA_7_SEGMENTE OF FPGA_7_SEGMENTE IS
signal refresh_counter: STD_LOGIC_VECTOR (19 downto 0);
signal LED_activating_counter: std_logic_vector(1 downto 0);
BEGIN
	process(clock)
	begin 
    if(CLOCK = '1' AND CLOCK'EVENT) then
        refresh_counter <= refresh_counter + 1;
    end if;
end process;
	LED_activating_counter <= refresh_counter(19 downto 18);
	process(LED_activating_counter)
begin
    case LED_activating_counter is
    when "00" =>
        Anode <= "0111"; 
        LED_OUT <= PRET_Z;
    when "01" =>
        Anode <= "1011"; 
        LED_OUT <= PRET_U;
    when "10" =>
        Anode <= "1101"; 
        LED_OUT <= SUMA_Z;
    when OTHERS =>
        Anode <= "1110"; 
        LED_OUT <= SUMA_U;   
    end case;
end process; 
END ARHITECTURA_FPGA_7_SEGMENTE;